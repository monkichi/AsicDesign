module lab2Cell();


//Instantiate the cell


endmodule
